// ED2platform.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module ED2platform (
		input  wire        clk_clk,               //            clk.clk
		output wire [2:0]  lcd_base_ctrl_export,  //  lcd_base_ctrl.export
		output wire [2:0]  lcd_cmd_export,        //        lcd_cmd.export
		inout  wire [15:0] lcd_data_export,       //       lcd_data.export
		output wire [15:0] pen_smp_period_export, // pen_smp_period.export
		input  wire        reset_reset_n,         //          reset.reset_n
		inout  wire        sd_card_b_SD_cmd,      //        sd_card.b_SD_cmd
		inout  wire        sd_card_b_SD_dat,      //               .b_SD_dat
		inout  wire        sd_card_b_SD_dat3,     //               .b_SD_dat3
		output wire        sd_card_o_SD_clock,    //               .o_SD_clock
		output wire [12:0] sdram_wire_addr,       //     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,         //               .ba
		output wire        sdram_wire_cas_n,      //               .cas_n
		output wire        sdram_wire_cke,        //               .cke
		output wire        sdram_wire_cs_n,       //               .cs_n
		inout  wire [31:0] sdram_wire_dq,         //               .dq
		output wire [3:0]  sdram_wire_dqm,        //               .dqm
		output wire        sdram_wire_ras_n,      //               .ras_n
		output wire        sdram_wire_we_n,       //               .we_n
		output wire [2:0]  touch_ctrl_export,     //     touch_ctrl.export
		input  wire [1:0]  touch_msg_export,      //      touch_msg.export
		input  wire        touch_pen_intr_export  // touch_pen_intr.export
	);

	wire  [31:0] cpu_data_master_readdata;                                                               // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                            // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                            // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                                                // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                             // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                                   // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                                          // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                                  // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                              // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                        // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                                     // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                                         // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                            // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                                   // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                                 // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                              // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect;  // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata;    // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest; // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address;     // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read;        // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	wire   [3:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable;  // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write;       // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	wire  [31:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata;   // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid0_control_slave_readdata;                                        // sysid0:readdata -> mm_interconnect_0:sysid0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid0_control_slave_address;                                         // mm_interconnect_0:sysid0_control_slave_address -> sysid0:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                         // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                      // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                      // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                          // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                             // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                       // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                            // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                        // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                  // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                                    // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                 // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                     // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                        // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                                  // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                               // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                       // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                                   // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_tftlcd_data_s1_chipselect;                                            // mm_interconnect_0:tftlcd_data_s1_chipselect -> tftlcd_data:chipselect
	wire  [31:0] mm_interconnect_0_tftlcd_data_s1_readdata;                                              // tftlcd_data:readdata -> mm_interconnect_0:tftlcd_data_s1_readdata
	wire   [1:0] mm_interconnect_0_tftlcd_data_s1_address;                                               // mm_interconnect_0:tftlcd_data_s1_address -> tftlcd_data:address
	wire         mm_interconnect_0_tftlcd_data_s1_write;                                                 // mm_interconnect_0:tftlcd_data_s1_write -> tftlcd_data:write_n
	wire  [31:0] mm_interconnect_0_tftlcd_data_s1_writedata;                                             // mm_interconnect_0:tftlcd_data_s1_writedata -> tftlcd_data:writedata
	wire         mm_interconnect_0_touch_pen_intr_s1_chipselect;                                         // mm_interconnect_0:touch_pen_intr_s1_chipselect -> touch_pen_intr:chipselect
	wire  [31:0] mm_interconnect_0_touch_pen_intr_s1_readdata;                                           // touch_pen_intr:readdata -> mm_interconnect_0:touch_pen_intr_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_pen_intr_s1_address;                                            // mm_interconnect_0:touch_pen_intr_s1_address -> touch_pen_intr:address
	wire         mm_interconnect_0_touch_pen_intr_s1_write;                                              // mm_interconnect_0:touch_pen_intr_s1_write -> touch_pen_intr:write_n
	wire  [31:0] mm_interconnect_0_touch_pen_intr_s1_writedata;                                          // mm_interconnect_0:touch_pen_intr_s1_writedata -> touch_pen_intr:writedata
	wire         mm_interconnect_0_tftlcd_cmd_s1_chipselect;                                             // mm_interconnect_0:tftlcd_cmd_s1_chipselect -> tftlcd_cmd:chipselect
	wire  [31:0] mm_interconnect_0_tftlcd_cmd_s1_readdata;                                               // tftlcd_cmd:readdata -> mm_interconnect_0:tftlcd_cmd_s1_readdata
	wire   [1:0] mm_interconnect_0_tftlcd_cmd_s1_address;                                                // mm_interconnect_0:tftlcd_cmd_s1_address -> tftlcd_cmd:address
	wire         mm_interconnect_0_tftlcd_cmd_s1_write;                                                  // mm_interconnect_0:tftlcd_cmd_s1_write -> tftlcd_cmd:write_n
	wire  [31:0] mm_interconnect_0_tftlcd_cmd_s1_writedata;                                              // mm_interconnect_0:tftlcd_cmd_s1_writedata -> tftlcd_cmd:writedata
	wire         mm_interconnect_0_tftlcd_base_ctrl_s1_chipselect;                                       // mm_interconnect_0:tftlcd_base_ctrl_s1_chipselect -> tftlcd_base_ctrl:chipselect
	wire  [31:0] mm_interconnect_0_tftlcd_base_ctrl_s1_readdata;                                         // tftlcd_base_ctrl:readdata -> mm_interconnect_0:tftlcd_base_ctrl_s1_readdata
	wire   [1:0] mm_interconnect_0_tftlcd_base_ctrl_s1_address;                                          // mm_interconnect_0:tftlcd_base_ctrl_s1_address -> tftlcd_base_ctrl:address
	wire         mm_interconnect_0_tftlcd_base_ctrl_s1_write;                                            // mm_interconnect_0:tftlcd_base_ctrl_s1_write -> tftlcd_base_ctrl:write_n
	wire  [31:0] mm_interconnect_0_tftlcd_base_ctrl_s1_writedata;                                        // mm_interconnect_0:tftlcd_base_ctrl_s1_writedata -> tftlcd_base_ctrl:writedata
	wire  [31:0] mm_interconnect_0_touch_msg_s1_readdata;                                                // touch_msg:readdata -> mm_interconnect_0:touch_msg_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_msg_s1_address;                                                 // mm_interconnect_0:touch_msg_s1_address -> touch_msg:address
	wire         mm_interconnect_0_touch_ctrl_s1_chipselect;                                             // mm_interconnect_0:touch_ctrl_s1_chipselect -> touch_ctrl:chipselect
	wire  [31:0] mm_interconnect_0_touch_ctrl_s1_readdata;                                               // touch_ctrl:readdata -> mm_interconnect_0:touch_ctrl_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_ctrl_s1_address;                                                // mm_interconnect_0:touch_ctrl_s1_address -> touch_ctrl:address
	wire         mm_interconnect_0_touch_ctrl_s1_write;                                                  // mm_interconnect_0:touch_ctrl_s1_write -> touch_ctrl:write_n
	wire  [31:0] mm_interconnect_0_touch_ctrl_s1_writedata;                                              // mm_interconnect_0:touch_ctrl_s1_writedata -> touch_ctrl:writedata
	wire         mm_interconnect_0_timer_1s_s1_chipselect;                                               // mm_interconnect_0:timer_1s_s1_chipselect -> timer_1s:chipselect
	wire  [15:0] mm_interconnect_0_timer_1s_s1_readdata;                                                 // timer_1s:readdata -> mm_interconnect_0:timer_1s_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1s_s1_address;                                                  // mm_interconnect_0:timer_1s_s1_address -> timer_1s:address
	wire         mm_interconnect_0_timer_1s_s1_write;                                                    // mm_interconnect_0:timer_1s_s1_write -> timer_1s:write_n
	wire  [15:0] mm_interconnect_0_timer_1s_s1_writedata;                                                // mm_interconnect_0:timer_1s_s1_writedata -> timer_1s:writedata
	wire         mm_interconnect_0_timer_scrollx_s1_chipselect;                                          // mm_interconnect_0:timer_scrollX_s1_chipselect -> timer_scrollX:chipselect
	wire  [15:0] mm_interconnect_0_timer_scrollx_s1_readdata;                                            // timer_scrollX:readdata -> mm_interconnect_0:timer_scrollX_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_scrollx_s1_address;                                             // mm_interconnect_0:timer_scrollX_s1_address -> timer_scrollX:address
	wire         mm_interconnect_0_timer_scrollx_s1_write;                                               // mm_interconnect_0:timer_scrollX_s1_write -> timer_scrollX:write_n
	wire  [15:0] mm_interconnect_0_timer_scrollx_s1_writedata;                                           // mm_interconnect_0:timer_scrollX_s1_writedata -> timer_scrollX:writedata
	wire         mm_interconnect_0_timer_touch_s1_chipselect;                                            // mm_interconnect_0:timer_touch_s1_chipselect -> timer_touch:chipselect
	wire  [15:0] mm_interconnect_0_timer_touch_s1_readdata;                                              // timer_touch:readdata -> mm_interconnect_0:timer_touch_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_touch_s1_address;                                               // mm_interconnect_0:timer_touch_s1_address -> timer_touch:address
	wire         mm_interconnect_0_timer_touch_s1_write;                                                 // mm_interconnect_0:timer_touch_s1_write -> timer_touch:write_n
	wire  [15:0] mm_interconnect_0_timer_touch_s1_writedata;                                             // mm_interconnect_0:timer_touch_s1_writedata -> timer_touch:writedata
	wire         mm_interconnect_0_pen_smp_speed_s1_chipselect;                                          // mm_interconnect_0:pen_smp_speed_s1_chipselect -> pen_smp_speed:chipselect
	wire  [31:0] mm_interconnect_0_pen_smp_speed_s1_readdata;                                            // pen_smp_speed:readdata -> mm_interconnect_0:pen_smp_speed_s1_readdata
	wire   [1:0] mm_interconnect_0_pen_smp_speed_s1_address;                                             // mm_interconnect_0:pen_smp_speed_s1_address -> pen_smp_speed:address
	wire         mm_interconnect_0_pen_smp_speed_s1_write;                                               // mm_interconnect_0:pen_smp_speed_s1_write -> pen_smp_speed:write_n
	wire  [31:0] mm_interconnect_0_pen_smp_speed_s1_writedata;                                           // mm_interconnect_0:pen_smp_speed_s1_writedata -> pen_smp_speed:writedata
	wire         irq_mapper_receiver0_irq;                                                               // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                               // timer_1s:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                               // timer_scrollX:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                               // timer_touch:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                               // touch_pen_intr:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                                                            // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                                         // rst_controller:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, pen_smp_speed:reset_n, rst_translator:in_reset, sdram:reset_n, sysid0:reset_n, tftlcd_base_ctrl:reset_n, tftlcd_cmd:reset_n, tftlcd_data:reset_n, timer_1s:reset_n, timer_scrollX:reset_n, timer_touch:reset_n, touch_ctrl:reset_n, touch_msg:reset_n, touch_pen_intr:reset_n]
	wire         rst_controller_reset_out_reset_req;                                                     // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                                          // cpu:debug_reset_request -> rst_controller:reset_in1

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (clk_clk),                                                                                //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                                        //               reset.reset_n
		.b_SD_cmd             (sd_card_b_SD_cmd),                                                                       //         conduit_end.export
		.b_SD_dat             (sd_card_b_SD_dat),                                                                       //                    .export
		.b_SD_dat3            (sd_card_b_SD_dat3),                                                                      //                    .export
		.o_SD_clock           (sd_card_o_SD_clock)                                                                      //                    .export
	);

	ED2platform_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	ED2platform_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	ED2platform_pen_smp_speed pen_smp_speed (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pen_smp_speed_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pen_smp_speed_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pen_smp_speed_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pen_smp_speed_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pen_smp_speed_s1_readdata),   //                    .readdata
		.out_port   (pen_smp_period_export)                          // external_connection.export
	);

	ED2platform_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	ED2platform_sysid0 sysid0 (
		.clock    (clk_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid0_control_slave_address)   //              .address
	);

	ED2platform_tftlcd_base_ctrl tftlcd_base_ctrl (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_tftlcd_base_ctrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tftlcd_base_ctrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tftlcd_base_ctrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tftlcd_base_ctrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tftlcd_base_ctrl_s1_readdata),   //                    .readdata
		.out_port   (lcd_base_ctrl_export)                              // external_connection.export
	);

	ED2platform_tftlcd_base_ctrl tftlcd_cmd (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_tftlcd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tftlcd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tftlcd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tftlcd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tftlcd_cmd_s1_readdata),   //                    .readdata
		.out_port   (lcd_cmd_export)                              // external_connection.export
	);

	ED2platform_tftlcd_data tftlcd_data (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_tftlcd_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tftlcd_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tftlcd_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tftlcd_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tftlcd_data_s1_readdata),   //                    .readdata
		.bidir_port (lcd_data_export)                              // external_connection.export
	);

	ED2platform_timer_1s timer_1s (
		.clk        (clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1s_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1s_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1s_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1s_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1s_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                  //   irq.irq
	);

	ED2platform_timer_scrollX timer_scrollx (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_timer_scrollx_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_scrollx_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_scrollx_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_scrollx_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_scrollx_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                       //   irq.irq
	);

	ED2platform_timer_scrollX timer_touch (
		.clk        (clk_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_timer_touch_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_touch_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_touch_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_touch_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_touch_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                     //   irq.irq
	);

	ED2platform_tftlcd_base_ctrl touch_ctrl (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_touch_ctrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_ctrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_ctrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_ctrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_ctrl_s1_readdata),   //                    .readdata
		.out_port   (touch_ctrl_export)                           // external_connection.export
	);

	ED2platform_touch_msg touch_msg (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_touch_msg_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touch_msg_s1_readdata), //                    .readdata
		.in_port  (touch_msg_export)                         // external_connection.export
	);

	ED2platform_touch_pen_intr touch_pen_intr (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_touch_pen_intr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_pen_intr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_pen_intr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_pen_intr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_pen_intr_s1_readdata),   //                    .readdata
		.in_port    (touch_pen_intr_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                        //                 irq.irq
	);

	ED2platform_mm_interconnect_0 mm_interconnect_0 (
		.clk_100_clk_clk                                                      (clk_clk),                                                                                //                                              clk_100_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset                                (rst_controller_reset_out_reset),                                                         //                          cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                              (cpu_data_master_address),                                                                //                                          cpu_data_master.address
		.cpu_data_master_waitrequest                                          (cpu_data_master_waitrequest),                                                            //                                                         .waitrequest
		.cpu_data_master_byteenable                                           (cpu_data_master_byteenable),                                                             //                                                         .byteenable
		.cpu_data_master_read                                                 (cpu_data_master_read),                                                                   //                                                         .read
		.cpu_data_master_readdata                                             (cpu_data_master_readdata),                                                               //                                                         .readdata
		.cpu_data_master_readdatavalid                                        (cpu_data_master_readdatavalid),                                                          //                                                         .readdatavalid
		.cpu_data_master_write                                                (cpu_data_master_write),                                                                  //                                                         .write
		.cpu_data_master_writedata                                            (cpu_data_master_writedata),                                                              //                                                         .writedata
		.cpu_data_master_debugaccess                                          (cpu_data_master_debugaccess),                                                            //                                                         .debugaccess
		.cpu_instruction_master_address                                       (cpu_instruction_master_address),                                                         //                                   cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                   (cpu_instruction_master_waitrequest),                                                     //                                                         .waitrequest
		.cpu_instruction_master_read                                          (cpu_instruction_master_read),                                                            //                                                         .read
		.cpu_instruction_master_readdata                                      (cpu_instruction_master_readdata),                                                        //                                                         .readdata
		.cpu_instruction_master_readdatavalid                                 (cpu_instruction_master_readdatavalid),                                                   //                                                         .readdatavalid
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                                                         .write
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                                                         .read
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                                                         .readdata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                                                         .writedata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                                                         .byteenable
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                                                         .waitrequest
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  //                                                         .chipselect
		.cpu_debug_mem_slave_address                                          (mm_interconnect_0_cpu_debug_mem_slave_address),                                          //                                      cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                            (mm_interconnect_0_cpu_debug_mem_slave_write),                                            //                                                         .write
		.cpu_debug_mem_slave_read                                             (mm_interconnect_0_cpu_debug_mem_slave_read),                                             //                                                         .read
		.cpu_debug_mem_slave_readdata                                         (mm_interconnect_0_cpu_debug_mem_slave_readdata),                                         //                                                         .readdata
		.cpu_debug_mem_slave_writedata                                        (mm_interconnect_0_cpu_debug_mem_slave_writedata),                                        //                                                         .writedata
		.cpu_debug_mem_slave_byteenable                                       (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                                       //                                                         .byteenable
		.cpu_debug_mem_slave_waitrequest                                      (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                                      //                                                         .waitrequest
		.cpu_debug_mem_slave_debugaccess                                      (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                                      //                                                         .debugaccess
		.jtag_uart_avalon_jtag_slave_address                                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                                  //                              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                                    //                                                         .write
		.jtag_uart_avalon_jtag_slave_read                                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                     //                                                         .read
		.jtag_uart_avalon_jtag_slave_readdata                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                                 //                                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                                //                                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                              //                                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                               //                                                         .chipselect
		.pen_smp_speed_s1_address                                             (mm_interconnect_0_pen_smp_speed_s1_address),                                             //                                         pen_smp_speed_s1.address
		.pen_smp_speed_s1_write                                               (mm_interconnect_0_pen_smp_speed_s1_write),                                               //                                                         .write
		.pen_smp_speed_s1_readdata                                            (mm_interconnect_0_pen_smp_speed_s1_readdata),                                            //                                                         .readdata
		.pen_smp_speed_s1_writedata                                           (mm_interconnect_0_pen_smp_speed_s1_writedata),                                           //                                                         .writedata
		.pen_smp_speed_s1_chipselect                                          (mm_interconnect_0_pen_smp_speed_s1_chipselect),                                          //                                                         .chipselect
		.sdram_s1_address                                                     (mm_interconnect_0_sdram_s1_address),                                                     //                                                 sdram_s1.address
		.sdram_s1_write                                                       (mm_interconnect_0_sdram_s1_write),                                                       //                                                         .write
		.sdram_s1_read                                                        (mm_interconnect_0_sdram_s1_read),                                                        //                                                         .read
		.sdram_s1_readdata                                                    (mm_interconnect_0_sdram_s1_readdata),                                                    //                                                         .readdata
		.sdram_s1_writedata                                                   (mm_interconnect_0_sdram_s1_writedata),                                                   //                                                         .writedata
		.sdram_s1_byteenable                                                  (mm_interconnect_0_sdram_s1_byteenable),                                                  //                                                         .byteenable
		.sdram_s1_readdatavalid                                               (mm_interconnect_0_sdram_s1_readdatavalid),                                               //                                                         .readdatavalid
		.sdram_s1_waitrequest                                                 (mm_interconnect_0_sdram_s1_waitrequest),                                                 //                                                         .waitrequest
		.sdram_s1_chipselect                                                  (mm_interconnect_0_sdram_s1_chipselect),                                                  //                                                         .chipselect
		.sysid0_control_slave_address                                         (mm_interconnect_0_sysid0_control_slave_address),                                         //                                     sysid0_control_slave.address
		.sysid0_control_slave_readdata                                        (mm_interconnect_0_sysid0_control_slave_readdata),                                        //                                                         .readdata
		.tftlcd_base_ctrl_s1_address                                          (mm_interconnect_0_tftlcd_base_ctrl_s1_address),                                          //                                      tftlcd_base_ctrl_s1.address
		.tftlcd_base_ctrl_s1_write                                            (mm_interconnect_0_tftlcd_base_ctrl_s1_write),                                            //                                                         .write
		.tftlcd_base_ctrl_s1_readdata                                         (mm_interconnect_0_tftlcd_base_ctrl_s1_readdata),                                         //                                                         .readdata
		.tftlcd_base_ctrl_s1_writedata                                        (mm_interconnect_0_tftlcd_base_ctrl_s1_writedata),                                        //                                                         .writedata
		.tftlcd_base_ctrl_s1_chipselect                                       (mm_interconnect_0_tftlcd_base_ctrl_s1_chipselect),                                       //                                                         .chipselect
		.tftlcd_cmd_s1_address                                                (mm_interconnect_0_tftlcd_cmd_s1_address),                                                //                                            tftlcd_cmd_s1.address
		.tftlcd_cmd_s1_write                                                  (mm_interconnect_0_tftlcd_cmd_s1_write),                                                  //                                                         .write
		.tftlcd_cmd_s1_readdata                                               (mm_interconnect_0_tftlcd_cmd_s1_readdata),                                               //                                                         .readdata
		.tftlcd_cmd_s1_writedata                                              (mm_interconnect_0_tftlcd_cmd_s1_writedata),                                              //                                                         .writedata
		.tftlcd_cmd_s1_chipselect                                             (mm_interconnect_0_tftlcd_cmd_s1_chipselect),                                             //                                                         .chipselect
		.tftlcd_data_s1_address                                               (mm_interconnect_0_tftlcd_data_s1_address),                                               //                                           tftlcd_data_s1.address
		.tftlcd_data_s1_write                                                 (mm_interconnect_0_tftlcd_data_s1_write),                                                 //                                                         .write
		.tftlcd_data_s1_readdata                                              (mm_interconnect_0_tftlcd_data_s1_readdata),                                              //                                                         .readdata
		.tftlcd_data_s1_writedata                                             (mm_interconnect_0_tftlcd_data_s1_writedata),                                             //                                                         .writedata
		.tftlcd_data_s1_chipselect                                            (mm_interconnect_0_tftlcd_data_s1_chipselect),                                            //                                                         .chipselect
		.timer_1s_s1_address                                                  (mm_interconnect_0_timer_1s_s1_address),                                                  //                                              timer_1s_s1.address
		.timer_1s_s1_write                                                    (mm_interconnect_0_timer_1s_s1_write),                                                    //                                                         .write
		.timer_1s_s1_readdata                                                 (mm_interconnect_0_timer_1s_s1_readdata),                                                 //                                                         .readdata
		.timer_1s_s1_writedata                                                (mm_interconnect_0_timer_1s_s1_writedata),                                                //                                                         .writedata
		.timer_1s_s1_chipselect                                               (mm_interconnect_0_timer_1s_s1_chipselect),                                               //                                                         .chipselect
		.timer_scrollX_s1_address                                             (mm_interconnect_0_timer_scrollx_s1_address),                                             //                                         timer_scrollX_s1.address
		.timer_scrollX_s1_write                                               (mm_interconnect_0_timer_scrollx_s1_write),                                               //                                                         .write
		.timer_scrollX_s1_readdata                                            (mm_interconnect_0_timer_scrollx_s1_readdata),                                            //                                                         .readdata
		.timer_scrollX_s1_writedata                                           (mm_interconnect_0_timer_scrollx_s1_writedata),                                           //                                                         .writedata
		.timer_scrollX_s1_chipselect                                          (mm_interconnect_0_timer_scrollx_s1_chipselect),                                          //                                                         .chipselect
		.timer_touch_s1_address                                               (mm_interconnect_0_timer_touch_s1_address),                                               //                                           timer_touch_s1.address
		.timer_touch_s1_write                                                 (mm_interconnect_0_timer_touch_s1_write),                                                 //                                                         .write
		.timer_touch_s1_readdata                                              (mm_interconnect_0_timer_touch_s1_readdata),                                              //                                                         .readdata
		.timer_touch_s1_writedata                                             (mm_interconnect_0_timer_touch_s1_writedata),                                             //                                                         .writedata
		.timer_touch_s1_chipselect                                            (mm_interconnect_0_timer_touch_s1_chipselect),                                            //                                                         .chipselect
		.touch_ctrl_s1_address                                                (mm_interconnect_0_touch_ctrl_s1_address),                                                //                                            touch_ctrl_s1.address
		.touch_ctrl_s1_write                                                  (mm_interconnect_0_touch_ctrl_s1_write),                                                  //                                                         .write
		.touch_ctrl_s1_readdata                                               (mm_interconnect_0_touch_ctrl_s1_readdata),                                               //                                                         .readdata
		.touch_ctrl_s1_writedata                                              (mm_interconnect_0_touch_ctrl_s1_writedata),                                              //                                                         .writedata
		.touch_ctrl_s1_chipselect                                             (mm_interconnect_0_touch_ctrl_s1_chipselect),                                             //                                                         .chipselect
		.touch_msg_s1_address                                                 (mm_interconnect_0_touch_msg_s1_address),                                                 //                                             touch_msg_s1.address
		.touch_msg_s1_readdata                                                (mm_interconnect_0_touch_msg_s1_readdata),                                                //                                                         .readdata
		.touch_pen_intr_s1_address                                            (mm_interconnect_0_touch_pen_intr_s1_address),                                            //                                        touch_pen_intr_s1.address
		.touch_pen_intr_s1_write                                              (mm_interconnect_0_touch_pen_intr_s1_write),                                              //                                                         .write
		.touch_pen_intr_s1_readdata                                           (mm_interconnect_0_touch_pen_intr_s1_readdata),                                           //                                                         .readdata
		.touch_pen_intr_s1_writedata                                          (mm_interconnect_0_touch_pen_intr_s1_writedata),                                          //                                                         .writedata
		.touch_pen_intr_s1_chipselect                                         (mm_interconnect_0_touch_pen_intr_s1_chipselect)                                          //                                                         .chipselect
	);

	ED2platform_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
